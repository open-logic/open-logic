Coverage Report Summary Data by instance

=================================================================================
=== Instance: /olo_base_cc_pulse_tb/i_dut/i_rst
=== Design Unit: olo.olo_base_cc_reset(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                        12        12         0   100.00%
    Statements                      12        12         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_pulse_tb/i_dut/i_sync/i_olo_base_cc_bits_constraints_region
=== Design Unit: olo.olo_base_cc_bits_constraints_entity(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       8         8         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_pulse_tb/i_dut
=== Design Unit: olo.olo_base_cc_pulse(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       9         9         0   100.00%

=================================================================================
=== Instance: /integer_vector_ptr_pkg
=== Design Unit: vunit_lib.integer_vector_ptr_pkg
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Assertions                       1         1         0   100.00%

=================================================================================
=== Instance: /string_ptr_pkg
=== Design Unit: vunit_lib.string_ptr_pkg
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Assertions                       1         1         0   100.00%

=================================================================================
=== Instance: /queue_pkg
=== Design Unit: vunit_lib.queue_pkg
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Assertions                       4         4         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_reset_tb/i_dut
=== Design Unit: olo.olo_base_cc_reset(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                        12        12         0   100.00%
    Statements                      12        12         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_status_tb/i_dut/i_scc/i_olo_base_cc_simple_constraints_region/i_pulse_cc/i_rst
=== Design Unit: olo.olo_base_cc_reset(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                        12        12         0   100.00%
    Statements                      12        12         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_status_tb/i_dut/i_scc/i_olo_base_cc_simple_constraints_region/i_pulse_cc/i_sync/i_olo_base_cc_bits_constraints_region
=== Design Unit: olo.olo_base_cc_bits_constraints_entity(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       8         8         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_status_tb/i_dut/i_scc/i_olo_base_cc_simple_constraints_region/i_pulse_cc
=== Design Unit: olo.olo_base_cc_pulse(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       9         9         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_status_tb/i_dut/i_scc/i_olo_base_cc_simple_constraints_region
=== Design Unit: olo.olo_base_cc_simple_constraints_entity(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         8         8         0   100.00%
    Statements                       7         7         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_status_tb/i_dut/i_bcc/i_rst
=== Design Unit: olo.olo_base_cc_reset(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                        12        12         0   100.00%
    Statements                      12        12         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_status_tb/i_dut/i_bcc/i_sync/i_olo_base_cc_bits_constraints_region
=== Design Unit: olo.olo_base_cc_bits_constraints_entity(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       8         8         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_status_tb/i_dut/i_bcc
=== Design Unit: olo.olo_base_cc_pulse(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       9         9         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_status_tb/i_dut
=== Design Unit: olo.olo_base_cc_status(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         5         5         0   100.00%
    Statements                       8         8         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_simple_tb/i_dut/i_olo_base_cc_simple_constraints_region/i_pulse_cc/i_rst
=== Design Unit: olo.olo_base_cc_reset(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                        12        12         0   100.00%
    Statements                      12        12         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_simple_tb/i_dut/i_olo_base_cc_simple_constraints_region/i_pulse_cc/i_sync/i_olo_base_cc_bits_constraints_region
=== Design Unit: olo.olo_base_cc_bits_constraints_entity(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       8         8         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_simple_tb/i_dut/i_olo_base_cc_simple_constraints_region/i_pulse_cc
=== Design Unit: olo.olo_base_cc_pulse(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       9         9         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_simple_tb/i_dut/i_olo_base_cc_simple_constraints_region
=== Design Unit: olo.olo_base_cc_simple_constraints_entity(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         8         8         0   100.00%
    Statements                       7         7         0   100.00%

=================================================================================
=== Instance: /olo_base_cc_bits_tb/i_dut/i_olo_base_cc_bits_constraints_region
=== Design Unit: olo.olo_base_cc_bits_constraints_entity(rtl)
=================================================================================
    Enabled Coverage              Bins      Hits    Misses  Coverage
    ----------------              ----      ----    ------  --------
    Branches                         6         6         0   100.00%
    Statements                       8         8         0   100.00%


TOTAL ASSERTION COVERAGE: 100.00%  ASSERTIONS: 6

Total Coverage By Instance (filtered view): 100.00%

