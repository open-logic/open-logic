---------------------------------------------------------------------------------------------------
-- Copyright (c) 2025 by Oliver Bründler
-- All rights reserved.
-- Authors: Milorad Petrovic
---------------------------------------------------------------------------------------------------

---------------------------------------------------------------------------------------------------
-- Libraries
---------------------------------------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

library vunit_lib;
    context vunit_lib.vunit_context;

library olo;
    use olo.olo_base_pkg_math.all;
    use olo.olo_base_pkg_logic.all;

---------------------------------------------------------------------------------------------------
-- Entity
---------------------------------------------------------------------------------------------------
entity olo_intf_inc_encoder_tb is
    generic (
        Clk_Frequency_g                : real                  := 100.0e6;
        DUT_PositionWidth_g            : natural               := 0;
        DUT_AngleWidth_g               : natural               := 0;
        EmulatedEncoder_ZPhaseExists_g : boolean               := FALSE;
        EmulatedEncoder_Resolution_g   : unsigned(63 downto 0);
        VUnit_WatchdogTimerDuration_g  : time                  := 10 ms;
        runner_cfg                     : string);
end entity;

architecture rtl of olo_intf_inc_encoder_tb is

    -- Main clock.
    constant Clk_Period_c : time := (1 sec) / Clk_Frequency_g;
    signal Clk : std_logic := '1';

    -- Phase signals generated by the emulated encoder.
    signal EmulatedEncoder_A : std_logic := '0';
    signal EmulatedEncoder_B : std_logic := '0';
    signal EmulatedEncoder_Z : std_logic := '0';

    -- Current angle of the emulated encoder.
    signal EmulatedEncoder_Angle : unsigned(EmulatedEncoder_Resolution_g'range) := (others => '0');

    -- DUT interface.
    signal DUT_Rst                  : std_logic := '1';
    signal DUT_Position_Value       : std_logic_vector(DUT_PositionWidth_g - 1 downto 0);
    signal DUT_Position_Clear       : std_logic := '0';
    signal DUT_Angle_Value          : std_logic_vector(DUT_AngleWidth_g - 1 downto 0);
    signal DUT_Angle_Clear          : std_logic := '0';
    signal DUT_Event_Up             : std_logic;
    signal DUT_Event_Down           : std_logic;
    signal DUT_Event_Index          : std_logic;

    -- This procedure waits for the specified number of clock rising edges.
    -- TODO: Move this procedure to the appropriate package.
    procedure WaitForClockCycles(
        signal   TargetClock               : in std_logic;
        constant NumberOfClockCyclesToWait : in positive) is
    begin

        -- Wait the requested number of clock cycles.
        for i in 1 to NumberOfClockCyclesToWait loop
            wait until rising_edge(TargetClock);
        end loop;

        -- There seems to be a bug in modelsim:
        -- The DUT outputs do not update instantaneously after a clock edge,
        -- hence this time wait is required so it is certain that all signals
        -- dependant on the clock edge are updated before any signal value checking is done.
        -- TODO: Further investigations of this issue are needed.
        wait for 1 ps;

    end procedure;

    -- This function calculates the remainded when dividing an numeric_std unsigned value
    -- with another numeric_std unsigned value. It is assumed that the dividend and divisor
    -- are of equal length, and a assert failure with occure if that is not provided.
    -- TODO: Move this procedure to the appropriate package.
    function UnsignedMod(
        Dividend : unsigned;
        Divisor  : unsigned
        ) return unsigned is
        variable Remainder : unsigned(Dividend'range) := Dividend;
    begin

        assert Dividend'length = Divisor'length report
            "Is is assumed that the dividend and divisor are of equal length."
            severity failure;

        while Remainder > Divisor loop
            Remainder := Remainder - Divisor;
        end loop;

        return Remainder;

    end function;

begin

    -- Instantiate VUnit watchdog timer.
    test_runner_watchdog(runner, VUnit_WatchdogTimerDuration_g);

    assert EmulatedEncoder_Resolution_g(1 downto 0) = "00" report
        "The value of the generic 'EmulatedEncoder_Resolution_g' is not valid. \n" &
        "The resolution of a quadrature encoder must be divisable by 4."
        severity error;

    proc_testcases : process is

        type EncoderStepDirection_t is (
            STEP_UP,
            STEP_DOWN);

        procedure RotateEncoder(
            StepDirection      : EncoderStepDirection_t;
            NumberOfSteps      : unsigned(63 downto 0) := to_unsigned(1, 64);
            ClockCyclesPerStep : positive := 1) is
            variable i : unsigned(63 downto 0);
        begin

            -- Rotate the encoder for the requested number of steps.
            i := NumberOfSteps;
            while i > 0 loop
                i := i - 1;

                if StepDirection = STEP_UP then
                    EmulatedEncoder_Angle <= (others => '0') when EmulatedEncoder_Angle = EmulatedEncoder_Resolution_g - 1 else EmulatedEncoder_Angle + 1;

                else -- StepDirection = STEP_DOWN
                    EmulatedEncoder_Angle <= EmulatedEncoder_Resolution_g - 1 when EmulatedEncoder_Angle = unsigned(zerosVector(EmulatedEncoder_Angle'length)) else EmulatedEncoder_Angle - 1;

                end if;

                WaitForClockCycles(Clk, ClockCyclesPerStep);

            end loop;

        end procedure;

        variable ExpectedAngleValue : unsigned(63 downto 0);

    begin
        test_runner_setup(runner, runner_cfg);

        set_stop_level(failure);

        while test_suite loop

            if run("ResetValues") then

                -- Check DUT outputs during reset.
                WaitForClockCycles(Clk, 1);
                check_equal(DUT_Position_Value, toUslv(0, DUT_PositionWidth_g), "DUT Position_Value is not zero during reset.");
                check_equal(DUT_Angle_Value, toUslv(0, DUT_AngleWidth_g), "DUT Angle_Value is not zero during reset.");
                check_equal(DUT_Event_Up, '0', "DUT Event_Up is not zero during reset.");
                check_equal(DUT_Event_Down, '0', "DUT Event_Down is not zero during reset.");
                check_equal(DUT_Event_Index, '0', "DUT Event_Index is not zero during reset.");

                -- Check DUT outputs right after releasing reset.
                DUT_Rst <= '0';
                WaitForClockCycles(Clk, 1);
                check_equal(DUT_Position_Value, toUslv(0, DUT_PositionWidth_g), "DUT Position_Value is not zero right after exiting reset.");
                check_equal(DUT_Angle_Value, toUslv(0, DUT_AngleWidth_g), "DUT Angle_Value is not zero right after exiting reset.");
                check_equal(DUT_Event_Up, '0', "DUT Event_Up is not zero right after exiting reset.");
                check_equal(DUT_Event_Down, '0', "DUT Event_Down is not zero right after exiting reset.");
                check_equal(DUT_Event_Index, '0', "DUT Event_Index is not zero right after exiting reset.");

            end if;

            if run("Basic") then

                -- Reset DUT, and then release reset.
                WaitForClockCycles(Clk, 1);
                DUT_Rst <= '0';

                -- Rotate encoder up for some amount.
                RotateEncoder(
                    StepDirection      => STEP_UP,
                    NumberOfSteps      => to_unsigned(10_000, 64),
                    ClockCyclesPerStep => 10);

                check_equal(DUT_Position_Value, toUslv(10_000, DUT_PositionWidth_g), "DUT 'Position_Value' is not the expected value after the positive direction rotation.");
                ExpectedAngleValue := UnsignedMod(to_unsigned(10_000, 64), EmulatedEncoder_Resolution_g);
                check_equal(DUT_Angle_Value, ExpectedAngleValue(DUT_Angle_Value'range), "DUT 'Angle_Value' is not the expected value after the positive direction rotation.");

                -- Rotate encoder down for some amount.
                RotateEncoder(
                    StepDirection      => STEP_DOWN,
                    NumberOfSteps      => to_unsigned(2_000, 64),
                    ClockCyclesPerStep => 10);

                check_equal(DUT_Position_Value, toUslv(8_000, DUT_PositionWidth_g), "DUT 'Position_Value' is not the expected value after the negative direction rotation.");
                ExpectedAngleValue := UnsignedMod(to_unsigned(8_000, 64), EmulatedEncoder_Resolution_g);
                check_equal(DUT_Angle_Value, ExpectedAngleValue(DUT_Angle_Value'range), "DUT 'Angle_Value' is not the expected value after the negative direction rotation.");

            end if;

            if run("EventGeneration") then

                -- Reset DUT, and then release reset.
                WaitForClockCycles(Clk, 1);
                DUT_Rst <= '0';

                -- Rotate in positive direction for some steps.
                for i in 1 to 10 loop
                    RotateEncoder(STEP_UP);
                    check_equal(DUT_Event_Up,    '1', "DUT did not signal an expected up count event.");
                    check_equal(DUT_Event_Down,  '0', "DUT signaled an unexpected down count event.");
                    check_equal(DUT_Event_Index, '0', "DUT signaled an unexpected index event.");
                    WaitForClockCycles(Clk, 9);
                end loop;

                -- Rotate in negative direction for some steps.
                for i in 1 to 5 loop
                    RotateEncoder(STEP_DOWN);
                    check_equal(DUT_Event_Up,    '0', "DUT signaled an unexpected up count event.");
                    check_equal(DUT_Event_Down,  '1', "DUT did not signal an expected down count event.");
                    check_equal(DUT_Event_Index, '0', "DUT signaled an unexpected index event.");
                    WaitForClockCycles(Clk, 9);
                end loop;

            end if;

            if run("AngleWrapAround") then

                -- Reset DUT, and then release reset.
                WaitForClockCycles(Clk, 1);
                DUT_Rst <= '0';

                -- Rotate up for a few steps.
                RotateEncoder(
                    StepDirection      => STEP_UP,
                    NumberOfSteps      => to_unsigned(10, 64),
                    ClockCyclesPerStep => 10);

                -- Rotate down just enough to wrap around.
                RotateEncoder(
                    StepDirection      => STEP_DOWN,
                    NumberOfSteps      => to_unsigned(11, 64),
                    ClockCyclesPerStep => 10);

                -- Check if angle value is as expected.
                check_equal(DUT_Angle_Value, resize(EmulatedEncoder_Resolution_g - 1, DUT_Angle_Value'length), "DUT angle value was not as expected.");

                -- Rotate down a little more.
                RotateEncoder(
                    StepDirection      => STEP_DOWN,
                    NumberOfSteps      => to_unsigned(5, 64),
                    ClockCyclesPerStep => 10);

                -- Rotate up just enough to wrap around.
                RotateEncoder(
                    StepDirection      => STEP_UP,
                    NumberOfSteps      => to_unsigned(6, 64),
                    ClockCyclesPerStep => 10);

                -- Check if angle value is as expected.
                check_equal(DUT_Angle_Value, to_unsigned(0, DUT_Angle_Value'length), "DUT angle value was not zero as expected.");

            end if;

            if run("AngleFullTurn") then

                -- Reset DUT, and then release reset.
                WaitForClockCycles(Clk, 1);
                DUT_Rst <= '0';

                -- Rotate up for one full turn.
                RotateEncoder(
                    StepDirection      => STEP_UP,
                    NumberOfSteps      => EmulatedEncoder_Resolution_g,
                    ClockCyclesPerStep => 10);

                -- DUT 'Angle_Value' should be zero.
                check_equal(DUT_Angle_Value, to_unsigned(0, DUT_Angle_Value'length), "DUT 'Angle_Value' was not zero as expected.");

                -- Rotate down for one full turn.
                RotateEncoder(
                    StepDirection      => STEP_DOWN,
                    NumberOfSteps      => EmulatedEncoder_Resolution_g,
                    ClockCyclesPerStep => 10);

                -- DUT 'Angle_Value' should be zero.
                check_equal(DUT_Angle_Value, to_unsigned(0, DUT_Angle_Value'length), "DUT 'Angle_Value' was not zero as expected.");

            end if;

        end loop;

        -- Wait for some idle cycles.
        WaitForClockCycles(Clk, 10);

        -- TB done
        test_runner_cleanup(runner);

    end process;

    -----------------------------------------------------------------------------------------------
    -- Clock
    -----------------------------------------------------------------------------------------------
    Clk <= not Clk after 0.5 * Clk_Period_c;

    -----------------------------------------------------------------------------------------------
    -- DUT
    -----------------------------------------------------------------------------------------------
    inst_dut : entity olo.olo_intf_inc_encoder
        generic map (
            AngleWidth_g    => DUT_AngleWidth_g,
            PositionWidth_g => DUT_PositionWidth_g)
        port map (
            Clk              => Clk,
            Rst              => DUT_Rst,
            Encoder_A        => EmulatedEncoder_A,
            Encoder_B        => EmulatedEncoder_B,
            Encoder_Z        => EmulatedEncoder_Z,
            Position_Value   => DUT_Position_Value,
            Position_Clear   => DUT_Position_Clear,
            Angle_Value      => DUT_Angle_Value,
            Angle_Clear      => DUT_Angle_Clear,
            Angle_Resolution => std_logic_vector(EmulatedEncoder_Resolution_g(DUT_AngleWidth_g downto 0)),
            Event_Up         => DUT_Event_Up,
            Event_Down       => DUT_Event_Down,
            Event_Index      => DUT_Event_Index
        );

    -----------------------------------------------------------------------------------------------
    -- Emulated encoder
    -----------------------------------------------------------------------------------------------
    proc_emulated_encoder : process (all) is
    begin

        -- Update encoder phases A and B.
        case EmulatedEncoder_Angle(1 downto 0) is

            when "00" =>
                EmulatedEncoder_A <= '0';
                EmulatedEncoder_B <= '0';

            when "01" =>
                EmulatedEncoder_A <= '1';
                EmulatedEncoder_B <= '0';

            when "10" =>
                EmulatedEncoder_A <= '1';
                EmulatedEncoder_B <= '1';

            when "11" =>
                EmulatedEncoder_A <= '0';
                EmulatedEncoder_B <= '1';

            when others =>
                check_failed("Emulated encoder angle is not a proper value!", failure);

        end case;

        -- Update encoder phase Z.
        EmulatedEncoder_Z <= '1' when EmulatedEncoder_ZPhaseExists_g and EmulatedEncoder_Angle = resize(EmulatedEncoder_Resolution_g - 1, EmulatedEncoder_Angle'length) else '0';

    end process;

end architecture rtl;
