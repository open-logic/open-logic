�      s`�,e F�e�8��&��tx��,���C#�80�3���%��'&Y&��X[Y�$ZX$[�&%3��d2  �L��   