---------------------------------------------------------------------------------------------------
-- Copyright (c) 2025 by Oliver Br�ndler, Switzerland
-- All rights reserved.
-- Authors: Oliver Bruendler
---------------------------------------------------------------------------------------------------

---------------------------------------------------------------------------------------------------
-- Libraries
---------------------------------------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

library vunit_lib;
    context vunit_lib.vunit_context;

library olo;
    use olo.olo_base_pkg_string.all;

---------------------------------------------------------------------------------------------------
-- Entity
---------------------------------------------------------------------------------------------------
-- vunit: run_all_in_same_sim
entity olo_base_pkg_string_tb is
    generic (
        runner_cfg     : string
    );
end entity;

architecture sim of olo_base_pkg_string_tb is

begin

    -----------------------------------------------------------------------------------------------
    -- TB Control
    -----------------------------------------------------------------------------------------------
    -- TB is not very vunit-ish because it is a package TB
    test_runner_watchdog(runner, 1 ms);

    p_control : process is
    begin
        test_runner_setup(runner, runner_cfg);

        wait for 1 ns;

        while test_suite loop

            if run("toUpper") then
                check_equal(toUpper("Hello"), "HELLO", "toUpper 1");
                check_equal(toUpper("hello"), "HELLO", "toUpper 2");
                check_equal(toUpper("hElLo"), "HELLO", "toUpper 3");
                check_equal(toUpper("HELLO"), "HELLO", "toUpper 4");
                check_equal(toUpper("123 &- abCD"), "123 ABCD", "toUpper 5");
            end if;

        end loop;

        wait for 1 ns;

        -- TB done
        test_runner_cleanup(runner);
    end process;

end architecture;
